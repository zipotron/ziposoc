module expander (input [16:0] instruction_C,
				 output [63:0] instruction);

endmodule
