module zipocpu (input clk,
				input [2:0] func,
				input sign,
				input [63:0] op_a,
				input [63:0] op_b,
				output reg [63:0] res);

endmodule
