flash_array[0]=32'h00000093;
flash_array[1]=32'h00000193;
flash_array[2]=32'h00000213;
flash_array[3]=32'h00000293;
flash_array[4]=32'h00000313;
flash_array[5]=32'h00000393;
flash_array[6]=32'h00000413;
flash_array[7]=32'h00000493;
flash_array[8]=32'h00000513;
flash_array[9]=32'h00000593;
flash_array[10]=32'h00000613;
flash_array[11]=32'h00000693;
flash_array[12]=32'h00000713;
flash_array[13]=32'h00000793;
flash_array[14]=32'h00000813;
flash_array[15]=32'h00000893;
flash_array[16]=32'h00000913;
flash_array[17]=32'h00000993;
flash_array[18]=32'h00000a13;
flash_array[19]=32'h00000a93;
flash_array[20]=32'h00000b13;
flash_array[21]=32'h00000b93;
flash_array[22]=32'h00000c13;
flash_array[23]=32'h00000c93;
flash_array[24]=32'h00000d13;
flash_array[25]=32'h00000d93;
flash_array[26]=32'h00000e13;
flash_array[27]=32'h00000e93;
flash_array[28]=32'h00000f13;
flash_array[29]=32'h00000f93;
flash_array[30]=32'h03000537;
flash_array[31]=32'hc10c4585;
flash_array[32]=32'hc1084501;
flash_array[33]=32'h4ee30511;
flash_array[34]=32'h0537fe25;
flash_array[35]=32'h458d0300;
flash_array[36]=32'h2011c10c;
flash_array[37]=32'h1101a001;
flash_array[38]=32'h1000ce22;
flash_array[39]=32'h030007b7;
flash_array[40]=32'h00078793;
flash_array[41]=32'hfef42223;
flash_array[42]=32'hfe042623;
flash_array[43]=32'h2783a819;
flash_array[44]=32'h0713fe44;
flash_array[45]=32'hc3980410;
flash_array[46]=32'hfec42783;
flash_array[47]=32'h26230785;
flash_array[48]=32'h2703fef4;
flash_array[49]=32'h6789fec4;
flash_array[50]=32'h70f78793;
flash_array[51]=32'hfee7d1e3;
flash_array[52]=32'hfe042423;
flash_array[53]=32'h2783a819;
flash_array[54]=32'h0713fe44;
flash_array[55]=32'hc3980810;
flash_array[56]=32'hfe842783;
flash_array[57]=32'h24230785;
flash_array[58]=32'h2703fef4;
flash_array[59]=32'h6789fe84;
flash_array[60]=32'h70f78793;
flash_array[61]=32'hfee7d1e3;
flash_array[62]=32'h0000bf45;
flash_array[63]=32'h00000000;
flash_array[64]=32'h00000000;
flash_array[65]=32'h00000000;
flash_array[66]=32'h00000000;
flash_array[67]=32'h00000000;
flash_array[68]=32'h00000000;
flash_array[69]=32'h00000000;
flash_array[70]=32'h00000000;
flash_array[71]=32'h00000000;
flash_array[72]=32'h00000000;
flash_array[73]=32'h00000000;
flash_array[74]=32'h00000000;
flash_array[75]=32'h00000000;
flash_array[76]=32'h00000000;
flash_array[77]=32'h00000000;
flash_array[78]=32'h00000000;
flash_array[79]=32'h00000000;
flash_array[80]=32'h00000000;
flash_array[81]=32'h00000000;
flash_array[82]=32'h00000000;
flash_array[83]=32'h00000000;
flash_array[84]=32'h00000000;
flash_array[85]=32'h00000000;
flash_array[86]=32'h00000000;
flash_array[87]=32'h00000000;
flash_array[88]=32'h00000000;
flash_array[89]=32'h00000000;
flash_array[90]=32'h00000000;
flash_array[91]=32'h00000000;
flash_array[92]=32'h00000000;
flash_array[93]=32'h00000000;
flash_array[94]=32'h00000000;
flash_array[95]=32'h00000000;
flash_array[96]=32'h00000000;
flash_array[97]=32'h00000000;
flash_array[98]=32'h00000000;
flash_array[99]=32'h00000000;
flash_array[100]=32'h00000000;
flash_array[101]=32'h00000000;
flash_array[102]=32'h00000000;
flash_array[103]=32'h00000000;
flash_array[104]=32'h00000000;
flash_array[105]=32'h00000000;
flash_array[106]=32'h00000000;
flash_array[107]=32'h00000000;
flash_array[108]=32'h00000000;
flash_array[109]=32'h00000000;
flash_array[110]=32'h00000000;
flash_array[111]=32'h00000000;
flash_array[112]=32'h00000000;
flash_array[113]=32'h00000000;
flash_array[114]=32'h00000000;
flash_array[115]=32'h00000000;
flash_array[116]=32'h00000000;
flash_array[117]=32'h00000000;
flash_array[118]=32'h00000000;
flash_array[119]=32'h00000000;
flash_array[120]=32'h00000000;
flash_array[121]=32'h00000000;
flash_array[122]=32'h00000000;
flash_array[123]=32'h00000000;
flash_array[124]=32'h00000000;
flash_array[125]=32'h00000000;
flash_array[126]=32'h00000000;
flash_array[127]=32'h00000000;
flash_array[128]=32'h00000000;
flash_array[129]=32'h00000000;
flash_array[130]=32'h00000000;
flash_array[131]=32'h00000000;
flash_array[132]=32'h00000000;
flash_array[133]=32'h00000000;
flash_array[134]=32'h00000000;
flash_array[135]=32'h00000000;
flash_array[136]=32'h00000000;
flash_array[137]=32'h00000000;
flash_array[138]=32'h00000000;
flash_array[139]=32'h00000000;
flash_array[140]=32'h00000000;
flash_array[141]=32'h00000000;
flash_array[142]=32'h00000000;
flash_array[143]=32'h00000000;
flash_array[144]=32'h00000000;
flash_array[145]=32'h00000000;
flash_array[146]=32'h00000000;
flash_array[147]=32'h00000000;
flash_array[148]=32'h00000000;
flash_array[149]=32'h00000000;
flash_array[150]=32'h00000000;
flash_array[151]=32'h00000000;
flash_array[152]=32'h00000000;
flash_array[153]=32'h00000000;
flash_array[154]=32'h00000000;
flash_array[155]=32'h00000000;
flash_array[156]=32'h00000000;
flash_array[157]=32'h00000000;
flash_array[158]=32'h00000000;
flash_array[159]=32'h00000000;
flash_array[160]=32'h00000000;
flash_array[161]=32'h00000000;
flash_array[162]=32'h00000000;
flash_array[163]=32'h00000000;
flash_array[164]=32'h00000000;
flash_array[165]=32'h00000000;
flash_array[166]=32'h00000000;
flash_array[167]=32'h00000000;
flash_array[168]=32'h00000000;
flash_array[169]=32'h00000000;
flash_array[170]=32'h00000000;
flash_array[171]=32'h00000000;
flash_array[172]=32'h00000000;
flash_array[173]=32'h00000000;
flash_array[174]=32'h00000000;
flash_array[175]=32'h00000000;
flash_array[176]=32'h00000000;
flash_array[177]=32'h00000000;
flash_array[178]=32'h00000000;
flash_array[179]=32'h00000000;
flash_array[180]=32'h00000000;
flash_array[181]=32'h00000000;
flash_array[182]=32'h00000000;
flash_array[183]=32'h00000000;
flash_array[184]=32'h00000000;
flash_array[185]=32'h00000000;
flash_array[186]=32'h00000000;
flash_array[187]=32'h00000000;
flash_array[188]=32'h00000000;
flash_array[189]=32'h00000000;
flash_array[190]=32'h00000000;
flash_array[191]=32'h00000000;
flash_array[192]=32'h00000000;
flash_array[193]=32'h00000000;
flash_array[194]=32'h00000000;
flash_array[195]=32'h00000000;
flash_array[196]=32'h00000000;
flash_array[197]=32'h00000000;
flash_array[198]=32'h00000000;
flash_array[199]=32'h00000000;
flash_array[200]=32'h00000000;
flash_array[201]=32'h00000000;
flash_array[202]=32'h00000000;
flash_array[203]=32'h00000000;
flash_array[204]=32'h00000000;
flash_array[205]=32'h00000000;
flash_array[206]=32'h00000000;
flash_array[207]=32'h00000000;
flash_array[208]=32'h00000000;
flash_array[209]=32'h00000000;
flash_array[210]=32'h00000000;
flash_array[211]=32'h00000000;
flash_array[212]=32'h00000000;
flash_array[213]=32'h00000000;
flash_array[214]=32'h00000000;
flash_array[215]=32'h00000000;
flash_array[216]=32'h00000000;
flash_array[217]=32'h00000000;
flash_array[218]=32'h00000000;
flash_array[219]=32'h00000000;
flash_array[220]=32'h00000000;
flash_array[221]=32'h00000000;
flash_array[222]=32'h00000000;
flash_array[223]=32'h00000000;
flash_array[224]=32'h00000000;
flash_array[225]=32'h00000000;
flash_array[226]=32'h00000000;
flash_array[227]=32'h00000000;
flash_array[228]=32'h00000000;
flash_array[229]=32'h00000000;
flash_array[230]=32'h00000000;
flash_array[231]=32'h00000000;
flash_array[232]=32'h00000000;
flash_array[233]=32'h00000000;
flash_array[234]=32'h00000000;
flash_array[235]=32'h00000000;
flash_array[236]=32'h00000000;
flash_array[237]=32'h00000000;
flash_array[238]=32'h00000000;
flash_array[239]=32'h00000000;
flash_array[240]=32'h00000000;
flash_array[241]=32'h00000000;
flash_array[242]=32'h00000000;
flash_array[243]=32'h00000000;
flash_array[244]=32'h00000000;
flash_array[245]=32'h00000000;
flash_array[246]=32'h00000000;
flash_array[247]=32'h00000000;
flash_array[248]=32'h00000000;
flash_array[249]=32'h00000000;
flash_array[250]=32'h00000000;
flash_array[251]=32'h00000000;
flash_array[252]=32'h00000000;
flash_array[253]=32'h00000000;
flash_array[254]=32'h00000000;
flash_array[255]=32'h00000000;
flash_array[256]=32'h00000000;
flash_array[257]=32'h00000000;
flash_array[258]=32'h00000000;
flash_array[259]=32'h00000000;
flash_array[260]=32'h00000000;
flash_array[261]=32'h00000000;
flash_array[262]=32'h00000000;
flash_array[263]=32'h00000000;
flash_array[264]=32'h00000000;
flash_array[265]=32'h00000000;
flash_array[266]=32'h00000000;
flash_array[267]=32'h00000000;
flash_array[268]=32'h00000000;
flash_array[269]=32'h00000000;
flash_array[270]=32'h00000000;
flash_array[271]=32'h00000000;
flash_array[272]=32'h00000000;
flash_array[273]=32'h00000000;
flash_array[274]=32'h00000000;
flash_array[275]=32'h00000000;
flash_array[276]=32'h00000000;
flash_array[277]=32'h00000000;
flash_array[278]=32'h00000000;
flash_array[279]=32'h00000000;
flash_array[280]=32'h00000000;
flash_array[281]=32'h00000000;
flash_array[282]=32'h00000000;
flash_array[283]=32'h00000000;
flash_array[284]=32'h00000000;
flash_array[285]=32'h00000000;
flash_array[286]=32'h00000000;
flash_array[287]=32'h00000000;
flash_array[288]=32'h00000000;
flash_array[289]=32'h00000000;
flash_array[290]=32'h00000000;
flash_array[291]=32'h00000000;
flash_array[292]=32'h00000000;
flash_array[293]=32'h00000000;
flash_array[294]=32'h00000000;
flash_array[295]=32'h00000000;
flash_array[296]=32'h00000000;
flash_array[297]=32'h00000000;
flash_array[298]=32'h00000000;
flash_array[299]=32'h00000000;
flash_array[300]=32'h00000000;
flash_array[301]=32'h00000000;
flash_array[302]=32'h00000000;
flash_array[303]=32'h00000000;
flash_array[304]=32'h00000000;
flash_array[305]=32'h00000000;
flash_array[306]=32'h00000000;
flash_array[307]=32'h00000000;
flash_array[308]=32'h00000000;
flash_array[309]=32'h00000000;
flash_array[310]=32'h00000000;
flash_array[311]=32'h00000000;
flash_array[312]=32'h00000000;
flash_array[313]=32'h00000000;
flash_array[314]=32'h00000000;
flash_array[315]=32'h00000000;
flash_array[316]=32'h00000000;
flash_array[317]=32'h00000000;
flash_array[318]=32'h00000000;
flash_array[319]=32'h00000000;
flash_array[320]=32'h00000000;
flash_array[321]=32'h00000000;
flash_array[322]=32'h00000000;
flash_array[323]=32'h00000000;
flash_array[324]=32'h00000000;
flash_array[325]=32'h00000000;
flash_array[326]=32'h00000000;
flash_array[327]=32'h00000000;
flash_array[328]=32'h00000000;
flash_array[329]=32'h00000000;
flash_array[330]=32'h00000000;
flash_array[331]=32'h00000000;
flash_array[332]=32'h00000000;
flash_array[333]=32'h00000000;
flash_array[334]=32'h00000000;
flash_array[335]=32'h00000000;
flash_array[336]=32'h00000000;
flash_array[337]=32'h00000000;
flash_array[338]=32'h00000000;
flash_array[339]=32'h00000000;
flash_array[340]=32'h00000000;
flash_array[341]=32'h00000000;
flash_array[342]=32'h00000000;
flash_array[343]=32'h00000000;
flash_array[344]=32'h00000000;
flash_array[345]=32'h00000000;
flash_array[346]=32'h00000000;
flash_array[347]=32'h00000000;
flash_array[348]=32'h00000000;
flash_array[349]=32'h00000000;
flash_array[350]=32'h00000000;
flash_array[351]=32'h00000000;
flash_array[352]=32'h00000000;
flash_array[353]=32'h00000000;
flash_array[354]=32'h00000000;
flash_array[355]=32'h00000000;
flash_array[356]=32'h00000000;
flash_array[357]=32'h00000000;
flash_array[358]=32'h00000000;
flash_array[359]=32'h00000000;
flash_array[360]=32'h00000000;
flash_array[361]=32'h00000000;
flash_array[362]=32'h00000000;
flash_array[363]=32'h00000000;
flash_array[364]=32'h00000000;
flash_array[365]=32'h00000000;
flash_array[366]=32'h00000000;
flash_array[367]=32'h00000000;
flash_array[368]=32'h00000000;
flash_array[369]=32'h00000000;
flash_array[370]=32'h00000000;
flash_array[371]=32'h00000000;
flash_array[372]=32'h00000000;
flash_array[373]=32'h00000000;
flash_array[374]=32'h00000000;
flash_array[375]=32'h00000000;
flash_array[376]=32'h00000000;
flash_array[377]=32'h00000000;
flash_array[378]=32'h00000000;
flash_array[379]=32'h00000000;
flash_array[380]=32'h00000000;
flash_array[381]=32'h00000000;
flash_array[382]=32'h00000000;
flash_array[383]=32'h00000000;
flash_array[384]=32'h00000000;
flash_array[385]=32'h00000000;
flash_array[386]=32'h00000000;
flash_array[387]=32'h00000000;
flash_array[388]=32'h00000000;
flash_array[389]=32'h00000000;
flash_array[390]=32'h00000000;
flash_array[391]=32'h00000000;
flash_array[392]=32'h00000000;
flash_array[393]=32'h00000000;
flash_array[394]=32'h00000000;
flash_array[395]=32'h00000000;
flash_array[396]=32'h00000000;
flash_array[397]=32'h00000000;
flash_array[398]=32'h00000000;
flash_array[399]=32'h00000000;
flash_array[400]=32'h00000000;
flash_array[401]=32'h00000000;
flash_array[402]=32'h00000000;
flash_array[403]=32'h00000000;
flash_array[404]=32'h00000000;
flash_array[405]=32'h00000000;
flash_array[406]=32'h00000000;
flash_array[407]=32'h00000000;
flash_array[408]=32'h00000000;
flash_array[409]=32'h00000000;
flash_array[410]=32'h00000000;
flash_array[411]=32'h00000000;
flash_array[412]=32'h00000000;
flash_array[413]=32'h00000000;
flash_array[414]=32'h00000000;
flash_array[415]=32'h00000000;
flash_array[416]=32'h00000000;
flash_array[417]=32'h00000000;
flash_array[418]=32'h00000000;
flash_array[419]=32'h00000000;
flash_array[420]=32'h00000000;
flash_array[421]=32'h00000000;
flash_array[422]=32'h00000000;
flash_array[423]=32'h00000000;
flash_array[424]=32'h00000000;
flash_array[425]=32'h00000000;
flash_array[426]=32'h00000000;
flash_array[427]=32'h00000000;
flash_array[428]=32'h00000000;
flash_array[429]=32'h00000000;
flash_array[430]=32'h00000000;
flash_array[431]=32'h00000000;
flash_array[432]=32'h00000000;
flash_array[433]=32'h00000000;
flash_array[434]=32'h00000000;
flash_array[435]=32'h00000000;
flash_array[436]=32'h00000000;
flash_array[437]=32'h00000000;
flash_array[438]=32'h00000000;
flash_array[439]=32'h00000000;
flash_array[440]=32'h00000000;
flash_array[441]=32'h00000000;
flash_array[442]=32'h00000000;
flash_array[443]=32'h00000000;
flash_array[444]=32'h00000000;
flash_array[445]=32'h00000000;
flash_array[446]=32'h00000000;
flash_array[447]=32'h00000000;
flash_array[448]=32'h00000000;
flash_array[449]=32'h00000000;
flash_array[450]=32'h00000000;
flash_array[451]=32'h00000000;
flash_array[452]=32'h00000000;
flash_array[453]=32'h00000000;
flash_array[454]=32'h00000000;
flash_array[455]=32'h00000000;
flash_array[456]=32'h00000000;
flash_array[457]=32'h00000000;
flash_array[458]=32'h00000000;
flash_array[459]=32'h00000000;
flash_array[460]=32'h00000000;
flash_array[461]=32'h00000000;
flash_array[462]=32'h00000000;
flash_array[463]=32'h00000000;
flash_array[464]=32'h00000000;
flash_array[465]=32'h00000000;
flash_array[466]=32'h00000000;
flash_array[467]=32'h00000000;
flash_array[468]=32'h00000000;
flash_array[469]=32'h00000000;
flash_array[470]=32'h00000000;
flash_array[471]=32'h00000000;
flash_array[472]=32'h00000000;
flash_array[473]=32'h00000000;
flash_array[474]=32'h00000000;
flash_array[475]=32'h00000000;
flash_array[476]=32'h00000000;
flash_array[477]=32'h00000000;
flash_array[478]=32'h00000000;
flash_array[479]=32'h00000000;
flash_array[480]=32'h00000000;
flash_array[481]=32'h00000000;
flash_array[482]=32'h00000000;
flash_array[483]=32'h00000000;
flash_array[484]=32'h00000000;
flash_array[485]=32'h00000000;
flash_array[486]=32'h00000000;
flash_array[487]=32'h00000000;
flash_array[488]=32'h00000000;
flash_array[489]=32'h00000000;
flash_array[490]=32'h00000000;
flash_array[491]=32'h00000000;
flash_array[492]=32'h00000000;
flash_array[493]=32'h00000000;
flash_array[494]=32'h00000000;
flash_array[495]=32'h00000000;
flash_array[496]=32'h00000000;
flash_array[497]=32'h00000000;
flash_array[498]=32'h00000000;
flash_array[499]=32'h00000000;
flash_array[500]=32'h00000000;
flash_array[501]=32'h00000000;
flash_array[502]=32'h00000000;
flash_array[503]=32'h00000000;
flash_array[504]=32'h00000000;
flash_array[505]=32'h00000000;
flash_array[506]=32'h00000000;
flash_array[507]=32'h00000000;
flash_array[508]=32'h00000000;
flash_array[509]=32'h00000000;
flash_array[510]=32'h00000000;
flash_array[511]=32'h00000000;
