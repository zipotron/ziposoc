{ram_array[64],ram_array[65],ram_array[66],ram_array[67]}=32'h00000093;
{ram_array[68],ram_array[69],ram_array[70],ram_array[71]}=32'h00000193;
{ram_array[72],ram_array[73],ram_array[74],ram_array[75]}=32'h00000213;
{ram_array[76],ram_array[77],ram_array[78],ram_array[79]}=32'h00000293;
{ram_array[80],ram_array[81],ram_array[82],ram_array[83]}=32'h00000313;
{ram_array[84],ram_array[85],ram_array[86],ram_array[87]}=32'h00000393;
{ram_array[88],ram_array[89],ram_array[90],ram_array[91]}=32'h00000413;
{ram_array[92],ram_array[93],ram_array[94],ram_array[95]}=32'h00000493;
{ram_array[96],ram_array[97],ram_array[98],ram_array[99]}=32'h00000513;
{ram_array[100],ram_array[101],ram_array[102],ram_array[103]}=32'h00000593;
{ram_array[104],ram_array[105],ram_array[106],ram_array[107]}=32'h00000613;
{ram_array[108],ram_array[109],ram_array[110],ram_array[111]}=32'h00000693;
{ram_array[112],ram_array[113],ram_array[114],ram_array[115]}=32'h00000713;
{ram_array[116],ram_array[117],ram_array[118],ram_array[119]}=32'h00000793;
{ram_array[120],ram_array[121],ram_array[122],ram_array[123]}=32'h00000813;
{ram_array[124],ram_array[125],ram_array[126],ram_array[127]}=32'h00000893;
{ram_array[128],ram_array[129],ram_array[130],ram_array[131]}=32'h00000913;
{ram_array[132],ram_array[133],ram_array[134],ram_array[135]}=32'h00000993;
{ram_array[136],ram_array[137],ram_array[138],ram_array[139]}=32'h00000a13;
{ram_array[140],ram_array[141],ram_array[142],ram_array[143]}=32'h00000a93;
{ram_array[144],ram_array[145],ram_array[146],ram_array[147]}=32'h00000b13;
{ram_array[148],ram_array[149],ram_array[150],ram_array[151]}=32'h00000b93;
{ram_array[152],ram_array[153],ram_array[154],ram_array[155]}=32'h00000c13;
{ram_array[156],ram_array[157],ram_array[158],ram_array[159]}=32'h00000c93;
{ram_array[160],ram_array[161],ram_array[162],ram_array[163]}=32'h00000d13;
{ram_array[164],ram_array[165],ram_array[166],ram_array[167]}=32'h00000d93;
{ram_array[168],ram_array[169],ram_array[170],ram_array[171]}=32'h00000e13;
{ram_array[172],ram_array[173],ram_array[174],ram_array[175]}=32'h00000e93;
{ram_array[176],ram_array[177],ram_array[178],ram_array[179]}=32'h00000f13;
{ram_array[180],ram_array[181],ram_array[182],ram_array[183]}=32'h00000f93;
{ram_array[184],ram_array[185],ram_array[186],ram_array[187]}=32'h03000537;
{ram_array[188],ram_array[189],ram_array[190],ram_array[191]}=32'hc10c4585;
{ram_array[192],ram_array[193],ram_array[194],ram_array[195]}=32'hc1084501;
{ram_array[196],ram_array[197],ram_array[198],ram_array[199]}=32'h4ee30511;
{ram_array[200],ram_array[201],ram_array[202],ram_array[203]}=32'h0537fe25;
{ram_array[204],ram_array[205],ram_array[206],ram_array[207]}=32'h458d0300;
{ram_array[208],ram_array[209],ram_array[210],ram_array[211]}=32'h2011c10c;
{ram_array[212],ram_array[213],ram_array[214],ram_array[215]}=32'h1101a001;
{ram_array[216],ram_array[217],ram_array[218],ram_array[219]}=32'h1000ce22;
{ram_array[220],ram_array[221],ram_array[222],ram_array[223]}=32'h030007b7;
{ram_array[224],ram_array[225],ram_array[226],ram_array[227]}=32'h00078793;
{ram_array[228],ram_array[229],ram_array[230],ram_array[231]}=32'hfef42223;
{ram_array[232],ram_array[233],ram_array[234],ram_array[235]}=32'hfe042623;
{ram_array[236],ram_array[237],ram_array[238],ram_array[239]}=32'h2783a819;
{ram_array[240],ram_array[241],ram_array[242],ram_array[243]}=32'h0713fe44;
{ram_array[244],ram_array[245],ram_array[246],ram_array[247]}=32'hc3980410;
{ram_array[248],ram_array[249],ram_array[250],ram_array[251]}=32'hfec42783;
{ram_array[252],ram_array[253],ram_array[254],ram_array[255]}=32'h26230785;
{ram_array[256],ram_array[257],ram_array[258],ram_array[259]}=32'h2703fef4;
{ram_array[260],ram_array[261],ram_array[262],ram_array[263]}=32'h6789fec4;
{ram_array[264],ram_array[265],ram_array[266],ram_array[267]}=32'h70f78793;
{ram_array[268],ram_array[269],ram_array[270],ram_array[271]}=32'hfee7d1e3;
{ram_array[272],ram_array[273],ram_array[274],ram_array[275]}=32'hfe042423;
{ram_array[276],ram_array[277],ram_array[278],ram_array[279]}=32'h2783a819;
{ram_array[280],ram_array[281],ram_array[282],ram_array[283]}=32'h0713fe44;
{ram_array[284],ram_array[285],ram_array[286],ram_array[287]}=32'hc3980810;
{ram_array[288],ram_array[289],ram_array[290],ram_array[291]}=32'hfe842783;
{ram_array[292],ram_array[293],ram_array[294],ram_array[295]}=32'h24230785;
{ram_array[296],ram_array[297],ram_array[298],ram_array[299]}=32'h2703fef4;
{ram_array[300],ram_array[301],ram_array[302],ram_array[303]}=32'h6789fe84;
{ram_array[304],ram_array[305],ram_array[306],ram_array[307]}=32'h70f78793;
{ram_array[308],ram_array[309],ram_array[310],ram_array[311]}=32'hfee7d1e3;
{ram_array[312],ram_array[313],ram_array[314],ram_array[315]}=32'h0000bf45;
{ram_array[316],ram_array[317],ram_array[318],ram_array[319]}=32'h00000000;
{ram_array[320],ram_array[321],ram_array[322],ram_array[323]}=32'h00000000;
{ram_array[324],ram_array[325],ram_array[326],ram_array[327]}=32'h00000000;
{ram_array[328],ram_array[329],ram_array[330],ram_array[331]}=32'h00000000;
{ram_array[332],ram_array[333],ram_array[334],ram_array[335]}=32'h00000000;
{ram_array[336],ram_array[337],ram_array[338],ram_array[339]}=32'h00000000;
{ram_array[340],ram_array[341],ram_array[342],ram_array[343]}=32'h00000000;
{ram_array[344],ram_array[345],ram_array[346],ram_array[347]}=32'h00000000;
{ram_array[348],ram_array[349],ram_array[350],ram_array[351]}=32'h00000000;
{ram_array[352],ram_array[353],ram_array[354],ram_array[355]}=32'h00000000;
{ram_array[356],ram_array[357],ram_array[358],ram_array[359]}=32'h00000000;
{ram_array[360],ram_array[361],ram_array[362],ram_array[363]}=32'h00000000;
{ram_array[364],ram_array[365],ram_array[366],ram_array[367]}=32'h00000000;
{ram_array[368],ram_array[369],ram_array[370],ram_array[371]}=32'h00000000;
{ram_array[372],ram_array[373],ram_array[374],ram_array[375]}=32'h00000000;
{ram_array[376],ram_array[377],ram_array[378],ram_array[379]}=32'h00000000;
{ram_array[380],ram_array[381],ram_array[382],ram_array[383]}=32'h00000000;
{ram_array[384],ram_array[385],ram_array[386],ram_array[387]}=32'h00000000;
{ram_array[388],ram_array[389],ram_array[390],ram_array[391]}=32'h00000000;
{ram_array[392],ram_array[393],ram_array[394],ram_array[395]}=32'h00000000;
{ram_array[396],ram_array[397],ram_array[398],ram_array[399]}=32'h00000000;
{ram_array[400],ram_array[401],ram_array[402],ram_array[403]}=32'h00000000;
{ram_array[404],ram_array[405],ram_array[406],ram_array[407]}=32'h00000000;
{ram_array[408],ram_array[409],ram_array[410],ram_array[411]}=32'h00000000;
{ram_array[412],ram_array[413],ram_array[414],ram_array[415]}=32'h00000000;
{ram_array[416],ram_array[417],ram_array[418],ram_array[419]}=32'h00000000;
{ram_array[420],ram_array[421],ram_array[422],ram_array[423]}=32'h00000000;
{ram_array[424],ram_array[425],ram_array[426],ram_array[427]}=32'h00000000;
{ram_array[428],ram_array[429],ram_array[430],ram_array[431]}=32'h00000000;
{ram_array[432],ram_array[433],ram_array[434],ram_array[435]}=32'h00000000;
{ram_array[436],ram_array[437],ram_array[438],ram_array[439]}=32'h00000000;
{ram_array[440],ram_array[441],ram_array[442],ram_array[443]}=32'h00000000;
{ram_array[444],ram_array[445],ram_array[446],ram_array[447]}=32'h00000000;
{ram_array[448],ram_array[449],ram_array[450],ram_array[451]}=32'h00000000;
{ram_array[452],ram_array[453],ram_array[454],ram_array[455]}=32'h00000000;
{ram_array[456],ram_array[457],ram_array[458],ram_array[459]}=32'h00000000;
{ram_array[460],ram_array[461],ram_array[462],ram_array[463]}=32'h00000000;
{ram_array[464],ram_array[465],ram_array[466],ram_array[467]}=32'h00000000;
{ram_array[468],ram_array[469],ram_array[470],ram_array[471]}=32'h00000000;
{ram_array[472],ram_array[473],ram_array[474],ram_array[475]}=32'h00000000;
{ram_array[476],ram_array[477],ram_array[478],ram_array[479]}=32'h00000000;
{ram_array[480],ram_array[481],ram_array[482],ram_array[483]}=32'h00000000;
{ram_array[484],ram_array[485],ram_array[486],ram_array[487]}=32'h00000000;
{ram_array[488],ram_array[489],ram_array[490],ram_array[491]}=32'h00000000;
{ram_array[492],ram_array[493],ram_array[494],ram_array[495]}=32'h00000000;
{ram_array[496],ram_array[497],ram_array[498],ram_array[499]}=32'h00000000;
{ram_array[500],ram_array[501],ram_array[502],ram_array[503]}=32'h00000000;
{ram_array[504],ram_array[505],ram_array[506],ram_array[507]}=32'h00000000;
{ram_array[508],ram_array[509],ram_array[510],ram_array[511]}=32'h00000000;
{ram_array[512],ram_array[513],ram_array[514],ram_array[515]}=32'h00000000;
{ram_array[516],ram_array[517],ram_array[518],ram_array[519]}=32'h00000000;
{ram_array[520],ram_array[521],ram_array[522],ram_array[523]}=32'h00000000;
{ram_array[524],ram_array[525],ram_array[526],ram_array[527]}=32'h00000000;
{ram_array[528],ram_array[529],ram_array[530],ram_array[531]}=32'h00000000;
{ram_array[532],ram_array[533],ram_array[534],ram_array[535]}=32'h00000000;
{ram_array[536],ram_array[537],ram_array[538],ram_array[539]}=32'h00000000;
{ram_array[540],ram_array[541],ram_array[542],ram_array[543]}=32'h00000000;
{ram_array[544],ram_array[545],ram_array[546],ram_array[547]}=32'h00000000;
{ram_array[548],ram_array[549],ram_array[550],ram_array[551]}=32'h00000000;
{ram_array[552],ram_array[553],ram_array[554],ram_array[555]}=32'h00000000;
{ram_array[556],ram_array[557],ram_array[558],ram_array[559]}=32'h00000000;
{ram_array[560],ram_array[561],ram_array[562],ram_array[563]}=32'h00000000;
{ram_array[564],ram_array[565],ram_array[566],ram_array[567]}=32'h00000000;
{ram_array[568],ram_array[569],ram_array[570],ram_array[571]}=32'h00000000;
{ram_array[572],ram_array[573],ram_array[574],ram_array[575]}=32'h00000000;
{ram_array[576],ram_array[577],ram_array[578],ram_array[579]}=32'h00000000;
{ram_array[580],ram_array[581],ram_array[582],ram_array[583]}=32'h00000000;
{ram_array[584],ram_array[585],ram_array[586],ram_array[587]}=32'h00000000;
{ram_array[588],ram_array[589],ram_array[590],ram_array[591]}=32'h00000000;
{ram_array[592],ram_array[593],ram_array[594],ram_array[595]}=32'h00000000;
{ram_array[596],ram_array[597],ram_array[598],ram_array[599]}=32'h00000000;
{ram_array[600],ram_array[601],ram_array[602],ram_array[603]}=32'h00000000;
{ram_array[604],ram_array[605],ram_array[606],ram_array[607]}=32'h00000000;
{ram_array[608],ram_array[609],ram_array[610],ram_array[611]}=32'h00000000;
{ram_array[612],ram_array[613],ram_array[614],ram_array[615]}=32'h00000000;
{ram_array[616],ram_array[617],ram_array[618],ram_array[619]}=32'h00000000;
{ram_array[620],ram_array[621],ram_array[622],ram_array[623]}=32'h00000000;
{ram_array[624],ram_array[625],ram_array[626],ram_array[627]}=32'h00000000;
{ram_array[628],ram_array[629],ram_array[630],ram_array[631]}=32'h00000000;
{ram_array[632],ram_array[633],ram_array[634],ram_array[635]}=32'h00000000;
{ram_array[636],ram_array[637],ram_array[638],ram_array[639]}=32'h00000000;
{ram_array[640],ram_array[641],ram_array[642],ram_array[643]}=32'h00000000;
{ram_array[644],ram_array[645],ram_array[646],ram_array[647]}=32'h00000000;
{ram_array[648],ram_array[649],ram_array[650],ram_array[651]}=32'h00000000;
{ram_array[652],ram_array[653],ram_array[654],ram_array[655]}=32'h00000000;
{ram_array[656],ram_array[657],ram_array[658],ram_array[659]}=32'h00000000;
{ram_array[660],ram_array[661],ram_array[662],ram_array[663]}=32'h00000000;
{ram_array[664],ram_array[665],ram_array[666],ram_array[667]}=32'h00000000;
{ram_array[668],ram_array[669],ram_array[670],ram_array[671]}=32'h00000000;
{ram_array[672],ram_array[673],ram_array[674],ram_array[675]}=32'h00000000;
{ram_array[676],ram_array[677],ram_array[678],ram_array[679]}=32'h00000000;
{ram_array[680],ram_array[681],ram_array[682],ram_array[683]}=32'h00000000;
{ram_array[684],ram_array[685],ram_array[686],ram_array[687]}=32'h00000000;
{ram_array[688],ram_array[689],ram_array[690],ram_array[691]}=32'h00000000;
{ram_array[692],ram_array[693],ram_array[694],ram_array[695]}=32'h00000000;
{ram_array[696],ram_array[697],ram_array[698],ram_array[699]}=32'h00000000;
{ram_array[700],ram_array[701],ram_array[702],ram_array[703]}=32'h00000000;
{ram_array[704],ram_array[705],ram_array[706],ram_array[707]}=32'h00000000;
{ram_array[708],ram_array[709],ram_array[710],ram_array[711]}=32'h00000000;
{ram_array[712],ram_array[713],ram_array[714],ram_array[715]}=32'h00000000;
{ram_array[716],ram_array[717],ram_array[718],ram_array[719]}=32'h00000000;
{ram_array[720],ram_array[721],ram_array[722],ram_array[723]}=32'h00000000;
{ram_array[724],ram_array[725],ram_array[726],ram_array[727]}=32'h00000000;
{ram_array[728],ram_array[729],ram_array[730],ram_array[731]}=32'h00000000;
{ram_array[732],ram_array[733],ram_array[734],ram_array[735]}=32'h00000000;
{ram_array[736],ram_array[737],ram_array[738],ram_array[739]}=32'h00000000;
{ram_array[740],ram_array[741],ram_array[742],ram_array[743]}=32'h00000000;
{ram_array[744],ram_array[745],ram_array[746],ram_array[747]}=32'h00000000;
{ram_array[748],ram_array[749],ram_array[750],ram_array[751]}=32'h00000000;
{ram_array[752],ram_array[753],ram_array[754],ram_array[755]}=32'h00000000;
{ram_array[756],ram_array[757],ram_array[758],ram_array[759]}=32'h00000000;
{ram_array[760],ram_array[761],ram_array[762],ram_array[763]}=32'h00000000;
{ram_array[764],ram_array[765],ram_array[766],ram_array[767]}=32'h00000000;
{ram_array[768],ram_array[769],ram_array[770],ram_array[771]}=32'h00000000;
{ram_array[772],ram_array[773],ram_array[774],ram_array[775]}=32'h00000000;
{ram_array[776],ram_array[777],ram_array[778],ram_array[779]}=32'h00000000;
{ram_array[780],ram_array[781],ram_array[782],ram_array[783]}=32'h00000000;
{ram_array[784],ram_array[785],ram_array[786],ram_array[787]}=32'h00000000;
{ram_array[788],ram_array[789],ram_array[790],ram_array[791]}=32'h00000000;
{ram_array[792],ram_array[793],ram_array[794],ram_array[795]}=32'h00000000;
{ram_array[796],ram_array[797],ram_array[798],ram_array[799]}=32'h00000000;
{ram_array[800],ram_array[801],ram_array[802],ram_array[803]}=32'h00000000;
{ram_array[804],ram_array[805],ram_array[806],ram_array[807]}=32'h00000000;
{ram_array[808],ram_array[809],ram_array[810],ram_array[811]}=32'h00000000;
{ram_array[812],ram_array[813],ram_array[814],ram_array[815]}=32'h00000000;
{ram_array[816],ram_array[817],ram_array[818],ram_array[819]}=32'h00000000;
{ram_array[820],ram_array[821],ram_array[822],ram_array[823]}=32'h00000000;
{ram_array[824],ram_array[825],ram_array[826],ram_array[827]}=32'h00000000;
{ram_array[828],ram_array[829],ram_array[830],ram_array[831]}=32'h00000000;
{ram_array[832],ram_array[833],ram_array[834],ram_array[835]}=32'h00000000;
{ram_array[836],ram_array[837],ram_array[838],ram_array[839]}=32'h00000000;
{ram_array[840],ram_array[841],ram_array[842],ram_array[843]}=32'h00000000;
{ram_array[844],ram_array[845],ram_array[846],ram_array[847]}=32'h00000000;
{ram_array[848],ram_array[849],ram_array[850],ram_array[851]}=32'h00000000;
{ram_array[852],ram_array[853],ram_array[854],ram_array[855]}=32'h00000000;
{ram_array[856],ram_array[857],ram_array[858],ram_array[859]}=32'h00000000;
{ram_array[860],ram_array[861],ram_array[862],ram_array[863]}=32'h00000000;
{ram_array[864],ram_array[865],ram_array[866],ram_array[867]}=32'h00000000;
{ram_array[868],ram_array[869],ram_array[870],ram_array[871]}=32'h00000000;
{ram_array[872],ram_array[873],ram_array[874],ram_array[875]}=32'h00000000;
{ram_array[876],ram_array[877],ram_array[878],ram_array[879]}=32'h00000000;
{ram_array[880],ram_array[881],ram_array[882],ram_array[883]}=32'h00000000;
{ram_array[884],ram_array[885],ram_array[886],ram_array[887]}=32'h00000000;
{ram_array[888],ram_array[889],ram_array[890],ram_array[891]}=32'h00000000;
{ram_array[892],ram_array[893],ram_array[894],ram_array[895]}=32'h00000000;
{ram_array[896],ram_array[897],ram_array[898],ram_array[899]}=32'h00000000;
{ram_array[900],ram_array[901],ram_array[902],ram_array[903]}=32'h00000000;
{ram_array[904],ram_array[905],ram_array[906],ram_array[907]}=32'h00000000;
{ram_array[908],ram_array[909],ram_array[910],ram_array[911]}=32'h00000000;
{ram_array[912],ram_array[913],ram_array[914],ram_array[915]}=32'h00000000;
{ram_array[916],ram_array[917],ram_array[918],ram_array[919]}=32'h00000000;
{ram_array[920],ram_array[921],ram_array[922],ram_array[923]}=32'h00000000;
{ram_array[924],ram_array[925],ram_array[926],ram_array[927]}=32'h00000000;
{ram_array[928],ram_array[929],ram_array[930],ram_array[931]}=32'h00000000;
{ram_array[932],ram_array[933],ram_array[934],ram_array[935]}=32'h00000000;
{ram_array[936],ram_array[937],ram_array[938],ram_array[939]}=32'h00000000;
{ram_array[940],ram_array[941],ram_array[942],ram_array[943]}=32'h00000000;
{ram_array[944],ram_array[945],ram_array[946],ram_array[947]}=32'h00000000;
{ram_array[948],ram_array[949],ram_array[950],ram_array[951]}=32'h00000000;
{ram_array[952],ram_array[953],ram_array[954],ram_array[955]}=32'h00000000;
{ram_array[956],ram_array[957],ram_array[958],ram_array[959]}=32'h00000000;
{ram_array[960],ram_array[961],ram_array[962],ram_array[963]}=32'h00000000;
{ram_array[964],ram_array[965],ram_array[966],ram_array[967]}=32'h00000000;
{ram_array[968],ram_array[969],ram_array[970],ram_array[971]}=32'h00000000;
{ram_array[972],ram_array[973],ram_array[974],ram_array[975]}=32'h00000000;
{ram_array[976],ram_array[977],ram_array[978],ram_array[979]}=32'h00000000;
{ram_array[980],ram_array[981],ram_array[982],ram_array[983]}=32'h00000000;
{ram_array[984],ram_array[985],ram_array[986],ram_array[987]}=32'h00000000;
{ram_array[988],ram_array[989],ram_array[990],ram_array[991]}=32'h00000000;
{ram_array[992],ram_array[993],ram_array[994],ram_array[995]}=32'h00000000;
{ram_array[996],ram_array[997],ram_array[998],ram_array[999]}=32'h00000000;
{ram_array[1000],ram_array[1001],ram_array[1002],ram_array[1003]}=32'h00000000;
{ram_array[1004],ram_array[1005],ram_array[1006],ram_array[1007]}=32'h00000000;
{ram_array[1008],ram_array[1009],ram_array[1010],ram_array[1011]}=32'h00000000;
{ram_array[1012],ram_array[1013],ram_array[1014],ram_array[1015]}=32'h00000000;
{ram_array[1016],ram_array[1017],ram_array[1018],ram_array[1019]}=32'h00000000;
{ram_array[1020],ram_array[1021],ram_array[1022],ram_array[1023]}=32'h00000000;
{ram_array[1024],ram_array[1025],ram_array[1026],ram_array[1027]}=32'h00000000;
{ram_array[1028],ram_array[1029],ram_array[1030],ram_array[1031]}=32'h00000000;
{ram_array[1032],ram_array[1033],ram_array[1034],ram_array[1035]}=32'h00000000;
{ram_array[1036],ram_array[1037],ram_array[1038],ram_array[1039]}=32'h00000000;
{ram_array[1040],ram_array[1041],ram_array[1042],ram_array[1043]}=32'h00000000;
{ram_array[1044],ram_array[1045],ram_array[1046],ram_array[1047]}=32'h00000000;
{ram_array[1048],ram_array[1049],ram_array[1050],ram_array[1051]}=32'h00000000;
{ram_array[1052],ram_array[1053],ram_array[1054],ram_array[1055]}=32'h00000000;
{ram_array[1056],ram_array[1057],ram_array[1058],ram_array[1059]}=32'h00000000;
{ram_array[1060],ram_array[1061],ram_array[1062],ram_array[1063]}=32'h00000000;
{ram_array[1064],ram_array[1065],ram_array[1066],ram_array[1067]}=32'h00000000;
{ram_array[1068],ram_array[1069],ram_array[1070],ram_array[1071]}=32'h00000000;
{ram_array[1072],ram_array[1073],ram_array[1074],ram_array[1075]}=32'h00000000;
{ram_array[1076],ram_array[1077],ram_array[1078],ram_array[1079]}=32'h00000000;
{ram_array[1080],ram_array[1081],ram_array[1082],ram_array[1083]}=32'h00000000;
{ram_array[1084],ram_array[1085],ram_array[1086],ram_array[1087]}=32'h00000000;
{ram_array[1088],ram_array[1089],ram_array[1090],ram_array[1091]}=32'h00000000;
{ram_array[1092],ram_array[1093],ram_array[1094],ram_array[1095]}=32'h00000000;
{ram_array[1096],ram_array[1097],ram_array[1098],ram_array[1099]}=32'h00000000;
{ram_array[1100],ram_array[1101],ram_array[1102],ram_array[1103]}=32'h00000000;
{ram_array[1104],ram_array[1105],ram_array[1106],ram_array[1107]}=32'h00000000;
{ram_array[1108],ram_array[1109],ram_array[1110],ram_array[1111]}=32'h00000000;
{ram_array[1112],ram_array[1113],ram_array[1114],ram_array[1115]}=32'h00000000;
{ram_array[1116],ram_array[1117],ram_array[1118],ram_array[1119]}=32'h00000000;
{ram_array[1120],ram_array[1121],ram_array[1122],ram_array[1123]}=32'h00000000;
{ram_array[1124],ram_array[1125],ram_array[1126],ram_array[1127]}=32'h00000000;
{ram_array[1128],ram_array[1129],ram_array[1130],ram_array[1131]}=32'h00000000;
{ram_array[1132],ram_array[1133],ram_array[1134],ram_array[1135]}=32'h00000000;
{ram_array[1136],ram_array[1137],ram_array[1138],ram_array[1139]}=32'h00000000;
{ram_array[1140],ram_array[1141],ram_array[1142],ram_array[1143]}=32'h00000000;
{ram_array[1144],ram_array[1145],ram_array[1146],ram_array[1147]}=32'h00000000;
{ram_array[1148],ram_array[1149],ram_array[1150],ram_array[1151]}=32'h00000000;
{ram_array[1152],ram_array[1153],ram_array[1154],ram_array[1155]}=32'h00000000;
{ram_array[1156],ram_array[1157],ram_array[1158],ram_array[1159]}=32'h00000000;
{ram_array[1160],ram_array[1161],ram_array[1162],ram_array[1163]}=32'h00000000;
{ram_array[1164],ram_array[1165],ram_array[1166],ram_array[1167]}=32'h00000000;
{ram_array[1168],ram_array[1169],ram_array[1170],ram_array[1171]}=32'h00000000;
{ram_array[1172],ram_array[1173],ram_array[1174],ram_array[1175]}=32'h00000000;
{ram_array[1176],ram_array[1177],ram_array[1178],ram_array[1179]}=32'h00000000;
{ram_array[1180],ram_array[1181],ram_array[1182],ram_array[1183]}=32'h00000000;
{ram_array[1184],ram_array[1185],ram_array[1186],ram_array[1187]}=32'h00000000;
{ram_array[1188],ram_array[1189],ram_array[1190],ram_array[1191]}=32'h00000000;
{ram_array[1192],ram_array[1193],ram_array[1194],ram_array[1195]}=32'h00000000;
{ram_array[1196],ram_array[1197],ram_array[1198],ram_array[1199]}=32'h00000000;
{ram_array[1200],ram_array[1201],ram_array[1202],ram_array[1203]}=32'h00000000;
{ram_array[1204],ram_array[1205],ram_array[1206],ram_array[1207]}=32'h00000000;
{ram_array[1208],ram_array[1209],ram_array[1210],ram_array[1211]}=32'h00000000;
{ram_array[1212],ram_array[1213],ram_array[1214],ram_array[1215]}=32'h00000000;
{ram_array[1216],ram_array[1217],ram_array[1218],ram_array[1219]}=32'h00000000;
{ram_array[1220],ram_array[1221],ram_array[1222],ram_array[1223]}=32'h00000000;
{ram_array[1224],ram_array[1225],ram_array[1226],ram_array[1227]}=32'h00000000;
{ram_array[1228],ram_array[1229],ram_array[1230],ram_array[1231]}=32'h00000000;
{ram_array[1232],ram_array[1233],ram_array[1234],ram_array[1235]}=32'h00000000;
{ram_array[1236],ram_array[1237],ram_array[1238],ram_array[1239]}=32'h00000000;
{ram_array[1240],ram_array[1241],ram_array[1242],ram_array[1243]}=32'h00000000;
{ram_array[1244],ram_array[1245],ram_array[1246],ram_array[1247]}=32'h00000000;
{ram_array[1248],ram_array[1249],ram_array[1250],ram_array[1251]}=32'h00000000;
{ram_array[1252],ram_array[1253],ram_array[1254],ram_array[1255]}=32'h00000000;
{ram_array[1256],ram_array[1257],ram_array[1258],ram_array[1259]}=32'h00000000;
{ram_array[1260],ram_array[1261],ram_array[1262],ram_array[1263]}=32'h00000000;
{ram_array[1264],ram_array[1265],ram_array[1266],ram_array[1267]}=32'h00000000;
{ram_array[1268],ram_array[1269],ram_array[1270],ram_array[1271]}=32'h00000000;
{ram_array[1272],ram_array[1273],ram_array[1274],ram_array[1275]}=32'h00000000;
{ram_array[1276],ram_array[1277],ram_array[1278],ram_array[1279]}=32'h00000000;
{ram_array[1280],ram_array[1281],ram_array[1282],ram_array[1283]}=32'h00000000;
{ram_array[1284],ram_array[1285],ram_array[1286],ram_array[1287]}=32'h00000000;
{ram_array[1288],ram_array[1289],ram_array[1290],ram_array[1291]}=32'h00000000;
{ram_array[1292],ram_array[1293],ram_array[1294],ram_array[1295]}=32'h00000000;
{ram_array[1296],ram_array[1297],ram_array[1298],ram_array[1299]}=32'h00000000;
{ram_array[1300],ram_array[1301],ram_array[1302],ram_array[1303]}=32'h00000000;
{ram_array[1304],ram_array[1305],ram_array[1306],ram_array[1307]}=32'h00000000;
{ram_array[1308],ram_array[1309],ram_array[1310],ram_array[1311]}=32'h00000000;
{ram_array[1312],ram_array[1313],ram_array[1314],ram_array[1315]}=32'h00000000;
{ram_array[1316],ram_array[1317],ram_array[1318],ram_array[1319]}=32'h00000000;
{ram_array[1320],ram_array[1321],ram_array[1322],ram_array[1323]}=32'h00000000;
{ram_array[1324],ram_array[1325],ram_array[1326],ram_array[1327]}=32'h00000000;
{ram_array[1328],ram_array[1329],ram_array[1330],ram_array[1331]}=32'h00000000;
{ram_array[1332],ram_array[1333],ram_array[1334],ram_array[1335]}=32'h00000000;
{ram_array[1336],ram_array[1337],ram_array[1338],ram_array[1339]}=32'h00000000;
{ram_array[1340],ram_array[1341],ram_array[1342],ram_array[1343]}=32'h00000000;
{ram_array[1344],ram_array[1345],ram_array[1346],ram_array[1347]}=32'h00000000;
{ram_array[1348],ram_array[1349],ram_array[1350],ram_array[1351]}=32'h00000000;
{ram_array[1352],ram_array[1353],ram_array[1354],ram_array[1355]}=32'h00000000;
{ram_array[1356],ram_array[1357],ram_array[1358],ram_array[1359]}=32'h00000000;
{ram_array[1360],ram_array[1361],ram_array[1362],ram_array[1363]}=32'h00000000;
{ram_array[1364],ram_array[1365],ram_array[1366],ram_array[1367]}=32'h00000000;
{ram_array[1368],ram_array[1369],ram_array[1370],ram_array[1371]}=32'h00000000;
{ram_array[1372],ram_array[1373],ram_array[1374],ram_array[1375]}=32'h00000000;
{ram_array[1376],ram_array[1377],ram_array[1378],ram_array[1379]}=32'h00000000;
{ram_array[1380],ram_array[1381],ram_array[1382],ram_array[1383]}=32'h00000000;
{ram_array[1384],ram_array[1385],ram_array[1386],ram_array[1387]}=32'h00000000;
{ram_array[1388],ram_array[1389],ram_array[1390],ram_array[1391]}=32'h00000000;
{ram_array[1392],ram_array[1393],ram_array[1394],ram_array[1395]}=32'h00000000;
{ram_array[1396],ram_array[1397],ram_array[1398],ram_array[1399]}=32'h00000000;
{ram_array[1400],ram_array[1401],ram_array[1402],ram_array[1403]}=32'h00000000;
{ram_array[1404],ram_array[1405],ram_array[1406],ram_array[1407]}=32'h00000000;
{ram_array[1408],ram_array[1409],ram_array[1410],ram_array[1411]}=32'h00000000;
{ram_array[1412],ram_array[1413],ram_array[1414],ram_array[1415]}=32'h00000000;
{ram_array[1416],ram_array[1417],ram_array[1418],ram_array[1419]}=32'h00000000;
{ram_array[1420],ram_array[1421],ram_array[1422],ram_array[1423]}=32'h00000000;
{ram_array[1424],ram_array[1425],ram_array[1426],ram_array[1427]}=32'h00000000;
{ram_array[1428],ram_array[1429],ram_array[1430],ram_array[1431]}=32'h00000000;
{ram_array[1432],ram_array[1433],ram_array[1434],ram_array[1435]}=32'h00000000;
{ram_array[1436],ram_array[1437],ram_array[1438],ram_array[1439]}=32'h00000000;
{ram_array[1440],ram_array[1441],ram_array[1442],ram_array[1443]}=32'h00000000;
{ram_array[1444],ram_array[1445],ram_array[1446],ram_array[1447]}=32'h00000000;
{ram_array[1448],ram_array[1449],ram_array[1450],ram_array[1451]}=32'h00000000;
{ram_array[1452],ram_array[1453],ram_array[1454],ram_array[1455]}=32'h00000000;
{ram_array[1456],ram_array[1457],ram_array[1458],ram_array[1459]}=32'h00000000;
{ram_array[1460],ram_array[1461],ram_array[1462],ram_array[1463]}=32'h00000000;
{ram_array[1464],ram_array[1465],ram_array[1466],ram_array[1467]}=32'h00000000;
{ram_array[1468],ram_array[1469],ram_array[1470],ram_array[1471]}=32'h00000000;
{ram_array[1472],ram_array[1473],ram_array[1474],ram_array[1475]}=32'h00000000;
{ram_array[1476],ram_array[1477],ram_array[1478],ram_array[1479]}=32'h00000000;
{ram_array[1480],ram_array[1481],ram_array[1482],ram_array[1483]}=32'h00000000;
{ram_array[1484],ram_array[1485],ram_array[1486],ram_array[1487]}=32'h00000000;
{ram_array[1488],ram_array[1489],ram_array[1490],ram_array[1491]}=32'h00000000;
{ram_array[1492],ram_array[1493],ram_array[1494],ram_array[1495]}=32'h00000000;
{ram_array[1496],ram_array[1497],ram_array[1498],ram_array[1499]}=32'h00000000;
{ram_array[1500],ram_array[1501],ram_array[1502],ram_array[1503]}=32'h00000000;
{ram_array[1504],ram_array[1505],ram_array[1506],ram_array[1507]}=32'h00000000;
{ram_array[1508],ram_array[1509],ram_array[1510],ram_array[1511]}=32'h00000000;
{ram_array[1512],ram_array[1513],ram_array[1514],ram_array[1515]}=32'h00000000;
{ram_array[1516],ram_array[1517],ram_array[1518],ram_array[1519]}=32'h00000000;
{ram_array[1520],ram_array[1521],ram_array[1522],ram_array[1523]}=32'h00000000;
{ram_array[1524],ram_array[1525],ram_array[1526],ram_array[1527]}=32'h00000000;
{ram_array[1528],ram_array[1529],ram_array[1530],ram_array[1531]}=32'h00000000;
{ram_array[1532],ram_array[1533],ram_array[1534],ram_array[1535]}=32'h00000000;
{ram_array[1536],ram_array[1537],ram_array[1538],ram_array[1539]}=32'h00000000;
{ram_array[1540],ram_array[1541],ram_array[1542],ram_array[1543]}=32'h00000000;
{ram_array[1544],ram_array[1545],ram_array[1546],ram_array[1547]}=32'h00000000;
{ram_array[1548],ram_array[1549],ram_array[1550],ram_array[1551]}=32'h00000000;
{ram_array[1552],ram_array[1553],ram_array[1554],ram_array[1555]}=32'h00000000;
{ram_array[1556],ram_array[1557],ram_array[1558],ram_array[1559]}=32'h00000000;
{ram_array[1560],ram_array[1561],ram_array[1562],ram_array[1563]}=32'h00000000;
{ram_array[1564],ram_array[1565],ram_array[1566],ram_array[1567]}=32'h00000000;
{ram_array[1568],ram_array[1569],ram_array[1570],ram_array[1571]}=32'h00000000;
{ram_array[1572],ram_array[1573],ram_array[1574],ram_array[1575]}=32'h00000000;
{ram_array[1576],ram_array[1577],ram_array[1578],ram_array[1579]}=32'h00000000;
{ram_array[1580],ram_array[1581],ram_array[1582],ram_array[1583]}=32'h00000000;
{ram_array[1584],ram_array[1585],ram_array[1586],ram_array[1587]}=32'h00000000;
{ram_array[1588],ram_array[1589],ram_array[1590],ram_array[1591]}=32'h00000000;
{ram_array[1592],ram_array[1593],ram_array[1594],ram_array[1595]}=32'h00000000;
{ram_array[1596],ram_array[1597],ram_array[1598],ram_array[1599]}=32'h00000000;
{ram_array[1600],ram_array[1601],ram_array[1602],ram_array[1603]}=32'h00000000;
{ram_array[1604],ram_array[1605],ram_array[1606],ram_array[1607]}=32'h00000000;
{ram_array[1608],ram_array[1609],ram_array[1610],ram_array[1611]}=32'h00000000;
{ram_array[1612],ram_array[1613],ram_array[1614],ram_array[1615]}=32'h00000000;
{ram_array[1616],ram_array[1617],ram_array[1618],ram_array[1619]}=32'h00000000;
{ram_array[1620],ram_array[1621],ram_array[1622],ram_array[1623]}=32'h00000000;
{ram_array[1624],ram_array[1625],ram_array[1626],ram_array[1627]}=32'h00000000;
{ram_array[1628],ram_array[1629],ram_array[1630],ram_array[1631]}=32'h00000000;
{ram_array[1632],ram_array[1633],ram_array[1634],ram_array[1635]}=32'h00000000;
{ram_array[1636],ram_array[1637],ram_array[1638],ram_array[1639]}=32'h00000000;
{ram_array[1640],ram_array[1641],ram_array[1642],ram_array[1643]}=32'h00000000;
{ram_array[1644],ram_array[1645],ram_array[1646],ram_array[1647]}=32'h00000000;
{ram_array[1648],ram_array[1649],ram_array[1650],ram_array[1651]}=32'h00000000;
{ram_array[1652],ram_array[1653],ram_array[1654],ram_array[1655]}=32'h00000000;
{ram_array[1656],ram_array[1657],ram_array[1658],ram_array[1659]}=32'h00000000;
{ram_array[1660],ram_array[1661],ram_array[1662],ram_array[1663]}=32'h00000000;
{ram_array[1664],ram_array[1665],ram_array[1666],ram_array[1667]}=32'h00000000;
{ram_array[1668],ram_array[1669],ram_array[1670],ram_array[1671]}=32'h00000000;
{ram_array[1672],ram_array[1673],ram_array[1674],ram_array[1675]}=32'h00000000;
{ram_array[1676],ram_array[1677],ram_array[1678],ram_array[1679]}=32'h00000000;
{ram_array[1680],ram_array[1681],ram_array[1682],ram_array[1683]}=32'h00000000;
{ram_array[1684],ram_array[1685],ram_array[1686],ram_array[1687]}=32'h00000000;
{ram_array[1688],ram_array[1689],ram_array[1690],ram_array[1691]}=32'h00000000;
{ram_array[1692],ram_array[1693],ram_array[1694],ram_array[1695]}=32'h00000000;
{ram_array[1696],ram_array[1697],ram_array[1698],ram_array[1699]}=32'h00000000;
{ram_array[1700],ram_array[1701],ram_array[1702],ram_array[1703]}=32'h00000000;
{ram_array[1704],ram_array[1705],ram_array[1706],ram_array[1707]}=32'h00000000;
{ram_array[1708],ram_array[1709],ram_array[1710],ram_array[1711]}=32'h00000000;
{ram_array[1712],ram_array[1713],ram_array[1714],ram_array[1715]}=32'h00000000;
{ram_array[1716],ram_array[1717],ram_array[1718],ram_array[1719]}=32'h00000000;
{ram_array[1720],ram_array[1721],ram_array[1722],ram_array[1723]}=32'h00000000;
{ram_array[1724],ram_array[1725],ram_array[1726],ram_array[1727]}=32'h00000000;
{ram_array[1728],ram_array[1729],ram_array[1730],ram_array[1731]}=32'h00000000;
{ram_array[1732],ram_array[1733],ram_array[1734],ram_array[1735]}=32'h00000000;
{ram_array[1736],ram_array[1737],ram_array[1738],ram_array[1739]}=32'h00000000;
{ram_array[1740],ram_array[1741],ram_array[1742],ram_array[1743]}=32'h00000000;
{ram_array[1744],ram_array[1745],ram_array[1746],ram_array[1747]}=32'h00000000;
{ram_array[1748],ram_array[1749],ram_array[1750],ram_array[1751]}=32'h00000000;
{ram_array[1752],ram_array[1753],ram_array[1754],ram_array[1755]}=32'h00000000;
{ram_array[1756],ram_array[1757],ram_array[1758],ram_array[1759]}=32'h00000000;
{ram_array[1760],ram_array[1761],ram_array[1762],ram_array[1763]}=32'h00000000;
{ram_array[1764],ram_array[1765],ram_array[1766],ram_array[1767]}=32'h00000000;
{ram_array[1768],ram_array[1769],ram_array[1770],ram_array[1771]}=32'h00000000;
{ram_array[1772],ram_array[1773],ram_array[1774],ram_array[1775]}=32'h00000000;
{ram_array[1776],ram_array[1777],ram_array[1778],ram_array[1779]}=32'h00000000;
{ram_array[1780],ram_array[1781],ram_array[1782],ram_array[1783]}=32'h00000000;
{ram_array[1784],ram_array[1785],ram_array[1786],ram_array[1787]}=32'h00000000;
{ram_array[1788],ram_array[1789],ram_array[1790],ram_array[1791]}=32'h00000000;
{ram_array[1792],ram_array[1793],ram_array[1794],ram_array[1795]}=32'h00000000;
{ram_array[1796],ram_array[1797],ram_array[1798],ram_array[1799]}=32'h00000000;
{ram_array[1800],ram_array[1801],ram_array[1802],ram_array[1803]}=32'h00000000;
{ram_array[1804],ram_array[1805],ram_array[1806],ram_array[1807]}=32'h00000000;
{ram_array[1808],ram_array[1809],ram_array[1810],ram_array[1811]}=32'h00000000;
{ram_array[1812],ram_array[1813],ram_array[1814],ram_array[1815]}=32'h00000000;
{ram_array[1816],ram_array[1817],ram_array[1818],ram_array[1819]}=32'h00000000;
{ram_array[1820],ram_array[1821],ram_array[1822],ram_array[1823]}=32'h00000000;
{ram_array[1824],ram_array[1825],ram_array[1826],ram_array[1827]}=32'h00000000;
{ram_array[1828],ram_array[1829],ram_array[1830],ram_array[1831]}=32'h00000000;
{ram_array[1832],ram_array[1833],ram_array[1834],ram_array[1835]}=32'h00000000;
{ram_array[1836],ram_array[1837],ram_array[1838],ram_array[1839]}=32'h00000000;
{ram_array[1840],ram_array[1841],ram_array[1842],ram_array[1843]}=32'h00000000;
{ram_array[1844],ram_array[1845],ram_array[1846],ram_array[1847]}=32'h00000000;
{ram_array[1848],ram_array[1849],ram_array[1850],ram_array[1851]}=32'h00000000;
{ram_array[1852],ram_array[1853],ram_array[1854],ram_array[1855]}=32'h00000000;
{ram_array[1856],ram_array[1857],ram_array[1858],ram_array[1859]}=32'h00000000;
{ram_array[1860],ram_array[1861],ram_array[1862],ram_array[1863]}=32'h00000000;
{ram_array[1864],ram_array[1865],ram_array[1866],ram_array[1867]}=32'h00000000;
{ram_array[1868],ram_array[1869],ram_array[1870],ram_array[1871]}=32'h00000000;
{ram_array[1872],ram_array[1873],ram_array[1874],ram_array[1875]}=32'h00000000;
{ram_array[1876],ram_array[1877],ram_array[1878],ram_array[1879]}=32'h00000000;
{ram_array[1880],ram_array[1881],ram_array[1882],ram_array[1883]}=32'h00000000;
{ram_array[1884],ram_array[1885],ram_array[1886],ram_array[1887]}=32'h00000000;
{ram_array[1888],ram_array[1889],ram_array[1890],ram_array[1891]}=32'h00000000;
{ram_array[1892],ram_array[1893],ram_array[1894],ram_array[1895]}=32'h00000000;
{ram_array[1896],ram_array[1897],ram_array[1898],ram_array[1899]}=32'h00000000;
{ram_array[1900],ram_array[1901],ram_array[1902],ram_array[1903]}=32'h00000000;
{ram_array[1904],ram_array[1905],ram_array[1906],ram_array[1907]}=32'h00000000;
{ram_array[1908],ram_array[1909],ram_array[1910],ram_array[1911]}=32'h00000000;
{ram_array[1912],ram_array[1913],ram_array[1914],ram_array[1915]}=32'h00000000;
{ram_array[1916],ram_array[1917],ram_array[1918],ram_array[1919]}=32'h00000000;
{ram_array[1920],ram_array[1921],ram_array[1922],ram_array[1923]}=32'h00000000;
{ram_array[1924],ram_array[1925],ram_array[1926],ram_array[1927]}=32'h00000000;
{ram_array[1928],ram_array[1929],ram_array[1930],ram_array[1931]}=32'h00000000;
{ram_array[1932],ram_array[1933],ram_array[1934],ram_array[1935]}=32'h00000000;
{ram_array[1936],ram_array[1937],ram_array[1938],ram_array[1939]}=32'h00000000;
{ram_array[1940],ram_array[1941],ram_array[1942],ram_array[1943]}=32'h00000000;
{ram_array[1944],ram_array[1945],ram_array[1946],ram_array[1947]}=32'h00000000;
{ram_array[1948],ram_array[1949],ram_array[1950],ram_array[1951]}=32'h00000000;
{ram_array[1952],ram_array[1953],ram_array[1954],ram_array[1955]}=32'h00000000;
{ram_array[1956],ram_array[1957],ram_array[1958],ram_array[1959]}=32'h00000000;
{ram_array[1960],ram_array[1961],ram_array[1962],ram_array[1963]}=32'h00000000;
{ram_array[1964],ram_array[1965],ram_array[1966],ram_array[1967]}=32'h00000000;
{ram_array[1968],ram_array[1969],ram_array[1970],ram_array[1971]}=32'h00000000;
{ram_array[1972],ram_array[1973],ram_array[1974],ram_array[1975]}=32'h00000000;
{ram_array[1976],ram_array[1977],ram_array[1978],ram_array[1979]}=32'h00000000;
{ram_array[1980],ram_array[1981],ram_array[1982],ram_array[1983]}=32'h00000000;
{ram_array[1984],ram_array[1985],ram_array[1986],ram_array[1987]}=32'h00000000;
{ram_array[1988],ram_array[1989],ram_array[1990],ram_array[1991]}=32'h00000000;
{ram_array[1992],ram_array[1993],ram_array[1994],ram_array[1995]}=32'h00000000;
{ram_array[1996],ram_array[1997],ram_array[1998],ram_array[1999]}=32'h00000000;
{ram_array[2000],ram_array[2001],ram_array[2002],ram_array[2003]}=32'h00000000;
{ram_array[2004],ram_array[2005],ram_array[2006],ram_array[2007]}=32'h00000000;
{ram_array[2008],ram_array[2009],ram_array[2010],ram_array[2011]}=32'h00000000;
{ram_array[2012],ram_array[2013],ram_array[2014],ram_array[2015]}=32'h00000000;
{ram_array[2016],ram_array[2017],ram_array[2018],ram_array[2019]}=32'h00000000;
{ram_array[2020],ram_array[2021],ram_array[2022],ram_array[2023]}=32'h00000000;
{ram_array[2024],ram_array[2025],ram_array[2026],ram_array[2027]}=32'h00000000;
{ram_array[2028],ram_array[2029],ram_array[2030],ram_array[2031]}=32'h00000000;
{ram_array[2032],ram_array[2033],ram_array[2034],ram_array[2035]}=32'h00000000;
{ram_array[2036],ram_array[2037],ram_array[2038],ram_array[2039]}=32'h00000000;
{ram_array[2040],ram_array[2041],ram_array[2042],ram_array[2043]}=32'h00000000;
{ram_array[2044],ram_array[2045],ram_array[2046],ram_array[2047]}=32'h00000000;
{ram_array[2048],ram_array[2049],ram_array[2050],ram_array[2051]}=32'h00000000;
{ram_array[2052],ram_array[2053],ram_array[2054],ram_array[2055]}=32'h00000000;
{ram_array[2056],ram_array[2057],ram_array[2058],ram_array[2059]}=32'h00000000;
{ram_array[2060],ram_array[2061],ram_array[2062],ram_array[2063]}=32'h00000000;
{ram_array[2064],ram_array[2065],ram_array[2066],ram_array[2067]}=32'h00000000;
{ram_array[2068],ram_array[2069],ram_array[2070],ram_array[2071]}=32'h00000000;
{ram_array[2072],ram_array[2073],ram_array[2074],ram_array[2075]}=32'h00000000;
{ram_array[2076],ram_array[2077],ram_array[2078],ram_array[2079]}=32'h00000000;
{ram_array[2080],ram_array[2081],ram_array[2082],ram_array[2083]}=32'h00000000;
{ram_array[2084],ram_array[2085],ram_array[2086],ram_array[2087]}=32'h00000000;
{ram_array[2088],ram_array[2089],ram_array[2090],ram_array[2091]}=32'h00000000;
{ram_array[2092],ram_array[2093],ram_array[2094],ram_array[2095]}=32'h00000000;
{ram_array[2096],ram_array[2097],ram_array[2098],ram_array[2099]}=32'h00000000;
{ram_array[2100],ram_array[2101],ram_array[2102],ram_array[2103]}=32'h00000000;
{ram_array[2104],ram_array[2105],ram_array[2106],ram_array[2107]}=32'h00000000;
{ram_array[2108],ram_array[2109],ram_array[2110],ram_array[2111]}=32'h00000000;
